-- ADD Rs, Rd
-- Rd <- Rs + Rd

--T3      Rd <= Rs + Rd   REGS_Read1 <= '1';
--                        REGS_Read2 <= '1';
--                        ALU_OP <= OP;
--                        Load_Status <= '1';
--                        REGS_Write <= '1';
--                        Clear <= '1';
